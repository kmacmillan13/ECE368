---------------------------------------------------
-- School:     University of Massachusetts Dartmouth
-- Department: Computer and Electrical Engineering
-- Engineer:   Emily DeBoer and Kayla MacMillan
-- 
-- Create Date:    SPRING 2015
-- Module Name:    StallConditionReg
-- Project Name:   UMD_RISC16
-- Target Devices: Spartan-3E
-- Tool versions:  Xilinx ISE 14.7
-- Description:    Control stalls
---------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE work.UMDRISC_pkg.ALL;
use work.all;

entity StallConditionReg is
    Port ( 
			  --Inputs
			  ifstall: out STD_LOGIC
			  --outputs
			  
			  );
			  
end StallConditionReg;

architecture Structural of StallConditionReg is

begin


end Structural;

